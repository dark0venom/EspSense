00000000  63 6f 6e 65 63 74 69 78  00 00 00 02 00 01 00 00  |conectix........|
00000010  00 00 00 00 00 00 02 00  01 23 45 67 2a 69 6d 67  |.........#Eg*img|
00000020  00 02 00 00 57 69 32 6b  00 00 00 00 00 fb 04 00  |....Wi2k........|
00000030  00 00 00 00 00 fb 04 00  00 02 ff 3f 00 00 00 03  |...........?....|
00000040  ff ff f5 b6 01 01 01 01  01 01 01 01 01 01 01 01  |................|
00000050  01 01 01 01 00 00 00 00  00 00 00 00 00 00 00 00  |................|
00000060  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00000200  63 78 73 70 61 72 73 65  ff ff ff ff ff ff ff ff  |cxsparse........|
00000210  00 00 00 00 00 00 06 00  00 01 00 00 00 00 00 08  |................|
00000220  00 20 00 00 ff ff f4 6f  00 00 00 00 00 00 00 00  |. .....o........|
00000230  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00000600  00 00 00 04 00 00 10 05  00 00 20 06 ff ff ff ff  |.......... .....|
00000610  ff ff ff ff ff ff ff ff  ff ff ff ff ff ff ff ff  |................|
*
00000a00  42 0a 42 0a 42 0a 42 0a  42 0a 42 0a 42 0a 42 0a  |B.B.B.B.B.B.B.B.|
*
00000bf0  42 0a 42 0a 42 0a 42 0a  42 0a 42 0a 42 0a 55 aa  |B.B.B.B.B.B.B.U.|
00000c00  94 c4 00 00 00 00 00 00  3f 00 01 00 00 00 00 00  |........?.......|
00000c10  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00000e00  42 0a 42 0a 42 0a 42 0a  42 0a 42 0a 42 0a 42 0a  |B.B.B.B.B.B.B.B.|
*
00002a00  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00008800  42 0a 42 0a 42 0a 42 0a  42 0a 42 0a 42 0a 42 0a  |B.B.B.B.B.B.B.B.|
*
00008a00  57 45 56 82 00 00 00 00  00 00 00 00 00 00 00 00  |WEV.............|
00008a10  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
00008a20  00 00 00 00 00 00 00 00  00 02 00 00 3f 00 00 00  |............?...|
00008a30  ff 00 00 00 01 00 00 00  c1 3e 00 00 c1 3e 00 00  |.........>...>..|
00008a40  00 00 00 00 00 00 00 00  10 0e 00 00 00 00 00 00  |................|
00008a50  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00008a80  00 00 00 00 57 45 56 82  1e 13 08 00 00 20 00 00  |....WEV...... ..|
00008a90  00 00 00 00 00 20 00 00  10 00 00 00 00 00 00 00  |..... ..........|
00008aa0  07 00 00 00 00 01 00 00  10 20 00 00 00 00 00 00  |......... ......|
00008ab0  01 00 00 00 c1 3e 00 00  00 00 00 00 00 00 00 00  |.....>..........|
00008ac0  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00008b10  00 00 00 00 42 0a 42 0a  42 0a 42 0a 42 0a 42 0a  |....B.B.B.B.B.B.|
00008b20  42 0a 42 0a 42 0a 42 0a  42 0a 42 0a 42 0a 42 0a  |B.B.B.B.B.B.B.B.|
*
0000a800  50 0a 50 0a 50 0a 50 0a  50 0a 50 0a 50 0a 50 0a  |P.P.P.P.P.P.P.P.|
*
00200a00  ff ff ff ff ff ff ff ff  ff ff ff ff ff ff ff ff  |................|
*
00200c00  50 0a 50 0a 50 0a 50 0a  50 0a 50 0a 50 0a 50 0a  |P.P.P.P.P.P.P.P.|
*
00400c00  ff ff ff ff ff ff ff ff  ff ff ff ff ff ff ff ff  |................|
*
00400e00  50 0a 50 0a 50 0a 50 0a  50 0a 50 0a 50 0a 50 0a  |P.P.P.P.P.P.P.P.|
*
0040ac00  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00650a00  63 6f 6e 65 63 74 69 78  00 00 00 02 00 01 00 00  |conectix........|
00650a10  00 00 00 00 00 00 02 00  01 23 45 67 2a 69 6d 67  |.........#Eg*img|
00650a20  00 02 00 00 57 69 32 6b  00 00 00 00 00 fb 04 00  |....Wi2k........|
00650a30  00 00 00 00 00 fb 04 00  00 02 ff 3f 00 00 00 03  |...........?....|
00650a40  ff ff f5 b6 01 01 01 01  01 01 01 01 01 01 01 01  |................|
00650a50  01 01 01 01 00 00 00 00  00 00 00 00 00 00 00 00  |................|
00650a60  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00650c00
