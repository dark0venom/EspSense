00000000  63 6f 6e 65 63 74 69 78  00 00 00 02 00 01 00 00  |conectix........|
00000010  00 00 00 00 00 00 02 00  01 23 45 67 2a 69 6d 67  |.........#Eg*img|
00000020  00 02 00 00 57 69 32 6b  00 00 00 00 00 7d 82 00  |....Wi2k.....}..|
00000030  00 00 00 00 00 7d 82 00  00 01 ff 3f 00 00 00 03  |.....}.....?....|
00000040  ff ff f5 87 04 04 04 04  04 04 04 04 04 04 04 04  |................|
00000050  04 04 04 04 00 00 00 00  00 00 00 00 00 00 00 00  |................|
00000060  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00000200  63 78 73 70 61 72 73 65  ff ff ff ff ff ff ff ff  |cxsparse........|
00000210  00 00 00 00 00 00 06 00  00 01 00 00 00 00 00 04  |................|
00000220  00 20 00 00 ff ff f4 73  00 00 00 00 00 00 00 00  |. .....s........|
00000230  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00000600  00 00 00 04 00 00 10 05  00 00 20 06 00 00 30 07  |.......... ...0.|
00000610  ff ff ff ff ff ff ff ff  ff ff ff ff ff ff ff ff  |................|
*
00000a00  42 0a 42 0a 42 0a 42 0a  42 0a 42 0a 42 0a 42 0a  |B.B.B.B.B.B.B.B.|
*
00000bb0  42 0a 42 0a 42 0a 42 0a  42 0a 42 0a 42 0a 00 00  |B.B.B.B.B.B.B...|
00000bc0  02 00 ee ff ff ff 01 00  00 00 c0 3e 00 00 00 00  |...........>....|
00000bd0  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00000bf0  00 00 00 00 00 00 00 00  00 00 00 00 00 00 55 aa  |..............U.|
00000c00  45 46 49 20 50 41 52 54  00 00 01 00 5c 00 00 00  |EFI PART....\...|
00000c10  0d 8a c6 7d 00 00 00 00  01 00 00 00 00 00 00 00  |...}............|
00000c20  c0 3e 00 00 00 00 00 00  03 00 00 00 00 00 00 00  |.>..............|
00000c30  be 3e 00 00 00 00 00 00  03 03 03 03 03 03 03 03  |.>..............|
00000c40  03 03 03 03 03 03 03 03  02 00 00 00 00 00 00 00  |................|
00000c50  02 00 00 00 80 00 00 00  3e b3 fa ad 00 00 00 00  |........>.......|
00000c60  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00000e00  b6 7c 6e 51 cf 6e d6 11  8f f8 00 02 2d 09 71 2b  |.|nQ.n......-.q+|
00000e10  01 01 01 01 01 01 01 01  01 01 01 01 01 01 01 01  |................|
00000e20  08 00 00 00 00 00 00 00  07 20 00 00 00 00 00 00  |......... ......|
00000e30  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00000e80  b5 7c 6e 51 cf 6e d6 11  8f f8 00 02 2d 09 71 2b  |.|nQ.n......-.q+|
00000e90  02 02 02 02 02 02 02 02  02 02 02 02 02 02 02 02  |................|
00000ea0  08 20 00 00 00 00 00 00  07 21 00 00 00 00 00 00  |. .......!......|
00000eb0  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00001a00  50 0a 50 0a 50 0a 50 0a  50 0a 50 0a 50 0a 50 0a  |P.P.P.P.P.P.P.P.|
*
00200a00  ff ff ff ff ff ff ff ff  ff ff ff ff ff ff ff ff  |................|
*
00200c00  50 0a 50 0a 50 0a 50 0a  50 0a 50 0a 50 0a 50 0a  |P.P.P.P.P.P.P.P.|
*
00400c00  ff ff ff ff ff ff ff ff  ff ff ff ff ff ff ff ff  |................|
*
00400e00  50 0a 50 0a 50 0a 50 0a  50 0a 50 0a 50 0a 50 0a  |P.P.P.P.P.P.P.P.|
*
00401e00  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00600e00  ff ff ff ff ff ff ff ff  ff ff ff ff ff ff ff ff  |................|
*
00601000  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
007d8e00  b6 7c 6e 51 cf 6e d6 11  8f f8 00 02 2d 09 71 2b  |.|nQ.n......-.q+|
007d8e10  01 01 01 01 01 01 01 01  01 01 01 01 01 01 01 01  |................|
007d8e20  08 00 00 00 00 00 00 00  07 20 00 00 00 00 00 00  |......... ......|
007d8e30  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
007d8e80  b5 7c 6e 51 cf 6e d6 11  8f f8 00 02 2d 09 71 2b  |.|nQ.n......-.q+|
007d8e90  02 02 02 02 02 02 02 02  02 02 02 02 02 02 02 02  |................|
007d8ea0  08 20 00 00 00 00 00 00  07 21 00 00 00 00 00 00  |. .......!......|
007d8eb0  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
007d9000  45 46 49 20 50 41 52 54  00 00 01 00 5c 00 00 00  |EFI PART....\...|
007d9010  19 14 f7 8a 00 00 00 00  c0 3e 00 00 00 00 00 00  |.........>......|
007d9020  01 00 00 00 00 00 00 00  03 00 00 00 00 00 00 00  |................|
007d9030  be 3e 00 00 00 00 00 00  03 03 03 03 03 03 03 03  |.>..............|
007d9040  03 03 03 03 03 03 03 03  bf 3e 00 00 00 00 00 00  |.........>......|
007d9050  02 00 00 00 80 00 00 00  3e b3 fa ad 00 00 00 00  |........>.......|
007d9060  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00801000  63 6f 6e 65 63 74 69 78  00 00 00 02 00 01 00 00  |conectix........|
00801010  00 00 00 00 00 00 02 00  01 23 45 67 2a 69 6d 67  |.........#Eg*img|
00801020  00 02 00 00 57 69 32 6b  00 00 00 00 00 7d 82 00  |....Wi2k.....}..|
00801030  00 00 00 00 00 7d 82 00  00 01 ff 3f 00 00 00 03  |.....}.....?....|
00801040  ff ff f5 87 04 04 04 04  04 04 04 04 04 04 04 04  |................|
00801050  04 04 04 04 00 00 00 00  00 00 00 00 00 00 00 00  |................|
00801060  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00801200
