00000000  63 6f 6e 65 63 74 69 78  00 00 00 02 00 01 00 00  |conectix........|
00000010  00 00 00 00 00 00 02 00  01 23 45 67 2a 69 6d 67  |.........#Eg*img|
00000020  00 02 00 00 57 69 32 6b  00 00 00 00 00 42 68 00  |....Wi2k.....Bh.|
00000030  00 00 00 00 00 42 68 00  00 7d 04 11 00 00 00 03  |.....Bh..}......|
00000040  ff ff f7 0e 01 01 01 01  01 01 01 01 01 01 01 01  |................|
00000050  01 01 01 01 00 00 00 00  00 00 00 00 00 00 00 00  |................|
00000060  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00000200  63 78 73 70 61 72 73 65  ff ff ff ff ff ff ff ff  |cxsparse........|
00000210  00 00 00 00 00 00 06 00  00 01 00 00 00 00 00 03  |................|
00000220  00 20 00 00 ff ff f4 74  00 00 00 00 00 00 00 00  |. .....t........|
00000230  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00000600  00 00 00 04 00 00 10 05  00 00 20 06 ff ff ff ff  |.......... .....|
00000610  ff ff ff ff ff ff ff ff  ff ff ff ff ff ff ff ff  |................|
*
00000a00  42 0a 42 0a 42 0a 42 0a  42 0a 42 0a 42 0a 42 0a  |B.B.B.B.B.B.B.B.|
*
00000bf0  42 0a 42 0a 42 0a 42 0a  42 0a 42 0a 42 0a 55 aa  |B.B.B.B.B.B.B.U.|
00000c00  94 c4 00 00 00 00 00 00  ff ff ff ff 00 00 00 00  |................|
00000c10  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00000e00  42 0a 42 0a 42 0a 42 0a  42 0a 42 0a 42 0a 42 0a  |B.B.B.B.B.B.B.B.|
*
00002c00  57 45 56 82 00 00 00 00  00 00 00 00 00 00 00 00  |WEV.............|
00002c10  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
00002c20  00 00 00 00 00 00 00 00  00 02 00 00 01 00 00 00  |................|
00002c30  01 00 00 00 10 21 00 00  01 00 00 00 10 21 00 00  |.....!.......!..|
00002c40  00 00 00 00 00 00 00 00  10 0e 00 00 00 00 00 00  |................|
00002c50  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00002c80  00 00 00 00 57 45 56 82  0f 0c 08 00 00 20 00 00  |....WEV...... ..|
00002c90  00 00 00 00 00 20 00 00  10 00 00 00 00 00 00 00  |..... ..........|
00002ca0  07 00 00 00 00 01 00 00  10 20 00 00 00 00 00 00  |......... ......|
00002cb0  01 00 00 00 10 21 00 00  00 00 00 00 00 00 00 00  |.....!..........|
00002cc0  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00002d10  00 00 00 00 42 0a 42 0a  42 0a 42 0a 42 0a 42 0a  |....B.B.B.B.B.B.|
00002d20  42 0a 42 0a 42 0a 42 0a  42 0a 42 0a 42 0a 42 0a  |B.B.B.B.B.B.B.B.|
*
00004a00  50 0a 50 0a 50 0a 50 0a  50 0a 50 0a 50 0a 50 0a  |P.P.P.P.P.P.P.P.|
*
00200a00  ff ff ff ff ff ff ff ff  ff ff ff ff ff ff ff ff  |................|
*
00200c00  50 0a 50 0a 50 0a 50 0a  50 0a 50 0a 50 0a 50 0a  |P.P.P.P.P.P.P.P.|
*
00400c00  ff ff ff ff ff ff ff ff  ff ff ff ff ff ff ff ff  |................|
*
00400e00  50 0a 50 0a 50 0a 50 0a  50 0a 50 0a 50 0a 50 0a  |P.P.P.P.P.P.P.P.|
*
00404e00  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00600e00  63 6f 6e 65 63 74 69 78  00 00 00 02 00 01 00 00  |conectix........|
00600e10  00 00 00 00 00 00 02 00  01 23 45 67 2a 69 6d 67  |.........#Eg*img|
00600e20  00 02 00 00 57 69 32 6b  00 00 00 00 00 42 68 00  |....Wi2k.....Bh.|
00600e30  00 00 00 00 00 42 68 00  00 7d 04 11 00 00 00 03  |.....Bh..}......|
00600e40  ff ff f7 0e 01 01 01 01  01 01 01 01 01 01 01 01  |................|
00600e50  01 01 01 01 00 00 00 00  00 00 00 00 00 00 00 00  |................|
00600e60  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00601000
