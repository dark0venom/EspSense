00000000  63 6f 6e 65 63 74 69 78  00 00 00 02 00 01 00 00  |conectix........|
00000010  00 00 00 00 00 00 02 00  01 23 45 67 2a 69 6d 67  |.........#Eg*img|
00000020  00 02 00 00 57 69 32 6b  00 00 00 00 00 42 68 00  |....Wi2k.....Bh.|
00000030  00 00 00 00 00 42 68 00  00 7d 04 11 00 00 00 03  |.....Bh..}......|
00000040  ff ff f6 de 04 04 04 04  04 04 04 04 04 04 04 04  |................|
00000050  04 04 04 04 00 00 00 00  00 00 00 00 00 00 00 00  |................|
00000060  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00000200  63 78 73 70 61 72 73 65  ff ff ff ff ff ff ff ff  |cxsparse........|
00000210  00 00 00 00 00 00 06 00  00 01 00 00 00 00 00 03  |................|
00000220  00 20 00 00 ff ff f4 74  00 00 00 00 00 00 00 00  |. .....t........|
00000230  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00000600  00 00 00 04 00 00 10 05  00 00 20 06 ff ff ff ff  |.......... .....|
00000610  ff ff ff ff ff ff ff ff  ff ff ff ff ff ff ff ff  |................|
*
00000a00  42 0a 42 0a 42 0a 42 0a  42 0a 42 0a 42 0a 42 0a  |B.B.B.B.B.B.B.B.|
*
00000bb0  42 0a 42 0a 42 0a 42 0a  42 0a 42 0a 42 0a 00 00  |B.B.B.B.B.B.B...|
00000bc0  02 00 ee ff ff ff 01 00  00 00 33 21 00 00 00 00  |..........3!....|
00000bd0  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00000bf0  00 00 00 00 00 00 00 00  00 00 00 00 00 00 55 aa  |..............U.|
00000c00  45 46 49 20 50 41 52 54  00 00 01 00 5c 00 00 00  |EFI PART....\...|
00000c10  c2 c7 92 19 00 00 00 00  01 00 00 00 00 00 00 00  |................|
00000c20  33 21 00 00 00 00 00 00  03 00 00 00 00 00 00 00  |3!..............|
00000c30  31 21 00 00 00 00 00 00  03 03 03 03 03 03 03 03  |1!..............|
00000c40  03 03 03 03 03 03 03 03  02 00 00 00 00 00 00 00  |................|
00000c50  02 00 00 00 80 00 00 00  3e b3 fa ad 00 00 00 00  |........>.......|
00000c60  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00000e00  b6 7c 6e 51 cf 6e d6 11  8f f8 00 02 2d 09 71 2b  |.|nQ.n......-.q+|
00000e10  01 01 01 01 01 01 01 01  01 01 01 01 01 01 01 01  |................|
00000e20  08 00 00 00 00 00 00 00  07 20 00 00 00 00 00 00  |......... ......|
00000e30  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00000e80  b5 7c 6e 51 cf 6e d6 11  8f f8 00 02 2d 09 71 2b  |.|nQ.n......-.q+|
00000e90  02 02 02 02 02 02 02 02  02 02 02 02 02 02 02 02  |................|
00000ea0  08 20 00 00 00 00 00 00  07 21 00 00 00 00 00 00  |. .......!......|
00000eb0  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00001a00  50 0a 50 0a 50 0a 50 0a  50 0a 50 0a 50 0a 50 0a  |P.P.P.P.P.P.P.P.|
*
00200a00  ff ff ff ff ff ff ff ff  ff ff ff ff ff ff ff ff  |................|
*
00200c00  50 0a 50 0a 50 0a 50 0a  50 0a 50 0a 50 0a 50 0a  |P.P.P.P.P.P.P.P.|
*
00400c00  ff ff ff ff ff ff ff ff  ff ff ff ff ff ff ff ff  |................|
*
00400e00  50 0a 50 0a 50 0a 50 0a  50 0a 50 0a 50 0a 50 0a  |P.P.P.P.P.P.P.P.|
*
00401e00  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00427200  b6 7c 6e 51 cf 6e d6 11  8f f8 00 02 2d 09 71 2b  |.|nQ.n......-.q+|
00427210  01 01 01 01 01 01 01 01  01 01 01 01 01 01 01 01  |................|
00427220  08 00 00 00 00 00 00 00  07 20 00 00 00 00 00 00  |......... ......|
00427230  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00427280  b5 7c 6e 51 cf 6e d6 11  8f f8 00 02 2d 09 71 2b  |.|nQ.n......-.q+|
00427290  02 02 02 02 02 02 02 02  02 02 02 02 02 02 02 02  |................|
004272a0  08 20 00 00 00 00 00 00  07 21 00 00 00 00 00 00  |. .......!......|
004272b0  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00427400  45 46 49 20 50 41 52 54  00 00 01 00 5c 00 00 00  |EFI PART....\...|
00427410  c0 86 13 46 00 00 00 00  33 21 00 00 00 00 00 00  |...F....3!......|
00427420  01 00 00 00 00 00 00 00  03 00 00 00 00 00 00 00  |................|
00427430  31 21 00 00 00 00 00 00  03 03 03 03 03 03 03 03  |1!..............|
00427440  03 03 03 03 03 03 03 03  32 21 00 00 00 00 00 00  |........2!......|
00427450  02 00 00 00 80 00 00 00  3e b3 fa ad 00 00 00 00  |........>.......|
00427460  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00600e00  63 6f 6e 65 63 74 69 78  00 00 00 02 00 01 00 00  |conectix........|
00600e10  00 00 00 00 00 00 02 00  01 23 45 67 2a 69 6d 67  |.........#Eg*img|
00600e20  00 02 00 00 57 69 32 6b  00 00 00 00 00 42 68 00  |....Wi2k.....Bh.|
00600e30  00 00 00 00 00 42 68 00  00 7d 04 11 00 00 00 03  |.....Bh..}......|
00600e40  ff ff f6 de 04 04 04 04  04 04 04 04 04 04 04 04  |................|
00600e50  04 04 04 04 00 00 00 00  00 00 00 00 00 00 00 00  |................|
00600e60  00 00 00 00 00 00 00 00  00 00 00 00 00 00 00 00  |................|
*
00601000
